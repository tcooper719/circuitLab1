module OR1 (output oor1, input A, B);
    assign oor1 = A | B;//this assigns the output oor1 to 
endmodule